lowConst_inst : lowConst PORT MAP (
		result	 => result_sig
	);
