constante_inst : constante PORT MAP (
		result	 => result_sig
	);
