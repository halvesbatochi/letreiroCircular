varedor_inst : varedor PORT MAP (
		clock	 => clock_sig,
		q	 => q_sig
	);
